module main(
    input clk_1hz,       // 1Hz ��ʱ�� (������ʱ��)
    input clk_1khz,      // 1000Hz ��Ƶʱ�� (���������ֵĽ���)
    input btn_1,     // Pulse 
    input btn_2,     // QD
    input btn_3_raw,     // CLR(��Ҫ��ת)
    input emergncy_stop, // ��ͣ����
    input switch_clr,      // ��λ����
    input simu_hopper_stop, // ©��ֹͣ�ź�
    input simu_hopper_add,  // ©���ֶ�����
    input simu_conveyor_stop, // ���ʹ�ֹͣ�ź�
    output [6:0] LED7S_out,
    output [3:0] LED7S2_out,
    output [3:0] LED7S3_out,
    output [3:0] LED7S4_out,
    output [3:0] LED7S5_out,
    output [3:0] LED7S6_out,
    output beep
);
    
    wire btn_3;
    assign btn_3 = ~btn_3_raw; // CLR����ȡ��������Ϊ�ߵ�ƽ

    // �򵥰��������ؼ�⣨ͬ���� clk_1khz��
    reg btn1_prev, btn2_prev;
    wire btn1_pressed = btn_1 && !btn1_prev;
    wire btn2_pressed = btn_2 && !btn2_prev;

    always @(posedge clk_1khz or negedge switch_clr) begin
        if (!switch_clr) begin
            btn1_prev <= 1'b0;
            btn2_prev <= 1'b0;
        end else begin
            btn1_prev <= btn_1;
            btn2_prev <= btn_2;
        end
    end

   
    // ==========================================
    // ��Ƶ
    // ==========================================
    reg [9:0] cnt1k;
    reg clk_4hz; // 4Hz ʱ�ӣ���������ܶ������������˸�ͷ�����
    reg clk_2hz; // 2Hz ʱ�ӣ���������ܷ�����
    reg clk_timer; // ��ʱ��ʱ�ӣ������л���ʱ����©����ʱ��

    always @(posedge clk_1khz) begin
        if (cnt1k == 1000-1) begin
            cnt1k <= 0;
            clk_timer <= ~clk_timer;
        end else
            cnt1k <= cnt1k + 1;
        
        if (cnt1k == 0 || cnt1k == 500)
            clk_2hz <= ~clk_2hz;
        
        if (cnt1k == 0 || cnt1k == 250 || cnt1k == 500 || cnt1k == 750)
            clk_4hz <= ~clk_4hz;
    end

    // ==========================================
    // ��״̬��
    // ==========================================
    
    reg [3:0] target_pills1; // �趨ÿƿҩƬ�� 0~999 ��λ
    reg [3:0] target_pills2; // �趨ÿƿҩƬ�� 0~999 ʮλ
    reg [3:0] target_pills3; // �趨ÿƿҩƬ�� 0~999 ��λ
    reg [3:0] target_bottles1; // �趨��ƿ�� 0~99 ��λ
    reg [3:0] target_bottles2; // �趨��ƿ�� 0~99 ʮλ
    reg [2:0] position; //��λ

    reg [3:0] now_pills1; // ��ǰƿҩƬ�� 0~999 ��λ
    reg [3:0] now_pills2; // ��ǰƿҩƬ�� 0~999 ʮλ
    reg [3:0] now_pills3; // ��ǰƿҩƬ�� 0~999 ��λ
    reg [3:0] now_bottles1; // �Ѿ���ɵ�ƿ�� 0~99 ��λ
    reg [3:0] now_bottles2; // �Ѿ���ɵ�ƿ�� 0~99 ʮλ

    // ״̬���壺�ϵ���� SETTING���� btn3 ȷ�Ͻ��� RUNNING���ﵽĿ��ƿ������ DONE
    localparam SETTING = 2'd0;
    localparam RUNNING = 2'd1;
    localparam DONE    = 2'd2;
    localparam ERROR   = 2'd3;

    reg [1:0] state;


    // Ŀ��/��ǰ��ֵ�Ա���ÿλ�Ĵ�����ʾ�������������ʾ��
    // ���Ƴ�©�������ؼ�⣨����ʱ��ʹ�ã�
    always @(posedge clk_1khz or negedge switch_clr) begin
        if (!switch_clr) begin
            state <= SETTING;
            // ���㵱ǰ����
            now_pills1 <= 4'd0; now_pills2 <= 4'd0; now_pills3 <= 4'd0;
            now_bottles1 <= 4'd0; now_bottles2 <= 4'd0;
            // ��ʼ��Ŀ��Ϊ
            target_pills1 <= 4'd1; target_pills2 <= 4'd0; target_pills3 <= 4'd0;
            target_bottles1 <= 4'd1; target_bottles2 <= 4'd0;
            position <= 3'd0;
        end else begin
            // ����̬��btn1 ��λ��btn2 ������ѡλ��btn3 ȷ�Ͽ�ʼ����
            if (state == SETTING) begin
                if (btn1_pressed) begin
                    // ѭ���л� 0..4��3λҩƬ + 2λƿ����
                    if (position == 3'd4) position <= 3'd0;
                    else position <= position + 1'b1;
                end

                if (btn2_pressed) begin
                    case (position)
                        3'd0: target_pills1 <= (target_pills1 == 4'd9) ? 4'd0 : target_pills1 + 1'b1;
                        3'd1: target_pills2 <= (target_pills2 == 4'd9) ? 4'd0 : target_pills2 + 1'b1;
                        3'd2: target_pills3 <= (target_pills3 == 4'd9) ? 4'd0 : target_pills3 + 1'b1;
                        3'd3: target_bottles1 <= (target_bottles1 == 4'd9) ? 4'd0 : target_bottles1 + 1'b1;
                        3'd4: target_bottles2 <= (target_bottles2 == 4'd9) ? 4'd0 : target_bottles2 + 1'b1;
                        default: ;
                    endcase
                end

                if (btn_3) begin
                    // ȷ�����ã��������ģʽ��RUNNING������ 0 ��ʼ����
                    state <= RUNNING;
                    now_pills1 <= 4'd0; now_pills2 <= 4'd0; now_pills3 <= 4'd0;
                    now_bottles1 <= 4'd0; now_bottles2 <= 4'd0;
                end
            end
            // ����̬��ȥ����©����ҩ�ͼ�ͣ�źŵ���������Ϊ�ֶ� btn2 ��Ϊ���Լ�������
            else if (state == RUNNING) begin
                // �����ã��� btn2 �ֶ�����ҩƬ������������֤�����߼���
                if (btn2_pressed) begin
                    // ����ҩƬ��������λ��λ��
                    if (now_pills1 == 4'd9) begin
                        now_pills1 <= 4'd0;
                        if (now_pills2 == 4'd9) begin
                            now_pills2 <= 4'd0;
                            if (now_pills3 == 4'd9) now_pills3 <= 4'd0;
                            else now_pills3 <= now_pills3 + 1'b1;
                        end else now_pills2 <= now_pills2 + 1'b1;
                    end else now_pills1 <= now_pills1 + 1'b1;

                    // �ж��Ƿ�ﵽĿ��ҩƬ�����Ƚ���λ��
                    if ((now_pills3 == target_pills3) && (now_pills2 == target_pills2) && (now_pills1 == target_pills1)) begin
                        // �ִ�Ŀ�꣺��ҩƬ����������ƿ������λ��λ��
                        now_pills1 <= 4'd0; now_pills2 <= 4'd0; now_pills3 <= 4'd0;
                        if (now_bottles1 == 4'd9) begin
                            now_bottles1 <= 4'd0;
                            now_bottles2 <= now_bottles2 + 1'b1;
                        end else now_bottles1 <= now_bottles1 + 1'b1;

                        // ����Ƿ�ﵽĿ��ƿ�����ﵽ����� DONE
                        if ((now_bottles2 == target_bottles2) && (now_bottles1 == target_bottles1)) begin
                            // �ﵽĿ��ƿ�� -> ���
                            state <= DONE;
                        end
                    end
                end

                
            end
            // ���̬���̰� btn3 ��������ģʽ�����õ�ǰ������
            else if (state == DONE) begin
                if (btn_3) begin
                    state <= SETTING;
                    now_pills1 <= 4'd0; now_pills2 <= 4'd0; now_pills3 <= 4'd0;
                    now_bottles1 <= 4'd0; now_bottles2 <= 4'd0;
                end
            end
            else if (state == ERROR) begin
                // ����̬���� btn3 ��������
                if (btn_3) begin
                    state <= SETTING;
                    now_pills1 <= 4'd0; now_pills2 <= 4'd0; now_pills3 <= 4'd0;
                    now_bottles1 <= 4'd0; now_bottles2 <= 4'd0;
                end
            end
        end
    end
    
    // ==========================================
    // ��ʾ����
    // ==========================================
    // �޸� display_1 ~ display_6 ��ֵ�����޸���ʾ����
    // �޸� flicker_mask[0...5] ��ֵ��������/�ر���˸


    wire [3:0] display_1;
    wire [3:0] display_2;
    wire [3:0] display_3;
    wire [3:0] display_4;
    wire [3:0] display_5;
    wire [3:0] display_6;

    // ������ʾ��SETTING ��ʾĿ�꣬����̬��ʾ��ǰ
    assign display_1 = state;
    assign display_2 = (state == SETTING) ? target_pills1   : now_pills1;
    assign display_3 = (state == SETTING) ? target_pills2   : now_pills2;
    assign display_4 = (state == SETTING) ? target_pills3   : now_pills3;
    assign display_5 = (state == SETTING) ? target_bottles1 : now_bottles1;
    assign display_6 = (state == SETTING) ? target_bottles2 : now_bottles2;

    reg [0:5] flicker_mask;

    assign LED7S2_out = (((~flicker_mask[1]) | clk_4hz) ? display_2 : 4'hf);
    assign LED7S3_out = (((~flicker_mask[2]) | clk_4hz) ? display_3 : 4'hf);
    assign LED7S4_out = (((~flicker_mask[3]) | clk_4hz) ? display_4 : 4'hf);
    assign LED7S5_out = (((~flicker_mask[4]) | clk_4hz) ? display_5 : 4'hf);
    assign LED7S6_out = (((~flicker_mask[5]) | clk_4hz) ? display_6 : 4'hf);
    assign LED7S_out = 7'b0000000;

    always @(*) begin
        if (state == SETTING) begin
            case (position)
                3'd0 : flicker_mask = 6'b010000;
                3'd1 : flicker_mask = 6'b001000;
                3'd2 : flicker_mask = 6'b000100;
                3'd3 : flicker_mask = 6'b000010;
                3'd4 : flicker_mask = 6'b000001;
            endcase
        end
        else begin
            flicker_mask = 6'b000000;
        end
            
    end
    // ==========================================
    // ���������֣��򻯣�DONE ʱ 2Hz ����������ʾ��
    // ==========================================
    // remove complex/undefined signals and keep simple behavior
    assign beep = (state == DONE) ? clk_2hz : 1'b0;

endmodule

