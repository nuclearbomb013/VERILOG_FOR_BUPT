module test(
    input clk,
    input clr,          // �ٶ�Ϊ�͵�ƽ��Ч (����ԭ���� negedge)
    output reg [6:0] LED7S,  // ����Ϊ��׼ [6:0] ��ʽ����λ�루�ֶ����룩
    output reg [3:0] LED7S2, // ʮλ�루BCD��
    output reg [3:0] LED7S3, // ��λ�֣�BCD��
    output reg [3:0] LED7S4, // ʮλ�֣�BCD��
    output reg [3:0] LED7S5, // ��λʱ��BCD��
    output reg [3:0] LED7S6  // ʮλʱ��BCD��
);

    reg [5:0] sec;
    reg [5:0] min;
    reg [4:0] hour;
    
    // ���ڸ����������ʱ����
    reg [3:0] sec_unit_val; 

    // ==========================================
    // 1. ʱ�Ӽ����븴λ�߼� (Clock and Reset)
    // ==========================================
    always @(posedge clk or negedge clr) begin
        if (!clr) begin
            // �첽��λ�����¸�λ��ʱ����
            sec <= 0;
            min <= 0;
            hour <= 0;
        end
        else begin
            // ���������߼�
            if (sec >= 59) begin
                sec <= 0;
                if (min >= 59) begin
                    min <= 0;
                    if (hour >= 23)
                        hour <= 0;
                    else
                        hour <= hour + 1;
                end
                else begin
                    min <= min + 1;
                end
            end
            else begin
                sec <= sec + 1;
            end
        end
    end

    // ==========================================
    // 2. ��λ����������߼� (Output Process)
    // ==========================================
    always @(*) begin
        // --- ��λ���벿�� (����������1) ---
        
        // �� (sec)
        sec_unit_val = sec % 10;     // ȡģ�ø�λ
        LED7S2       = sec / 10;     // ������ʮλ
        
        // �� (min)
        LED7S3       = min % 10;     // ��λ
        LED7S4       = min / 10;     // ʮλ
        
        // ʱ (hour)
        LED7S5       = hour % 10;    // ��λ
        LED7S6       = hour / 10;    // ʮλ

        // --- �ֶ����벿�� (�����ĸ�λ) ---
        // �����ǹ��������ǹ�����ȡ����Ӳ���������������ṩ�ı���
        // 4'b0000 -> 7'b1111110 (0x7E, �������������ĸߵ�ƽ�����������ǹ������ĵ͵�ƽ��Ч)
        case (sec_unit_val)
			4'd0: LED7S <= 7'b0111111; // 0: a,b,c,d,e,f ��
            4'd1: LED7S <= 7'b0000110; // 1: b,c ��
            4'd2: LED7S <= 7'b1011011; // 2: a,b,d,e,g ��
            4'd3: LED7S <= 7'b1001111; // 3: a,b,c,d,g ��
            4'd4: LED7S <= 7'b1100110; // 4: b,c,f,g ��
            4'd5: LED7S <= 7'b1101101; // 5: a,c,d,f,g ��
            4'd6: LED7S <= 7'b1111100; // 6: c,d,e,f,g ��
            4'd7: LED7S <= 7'b0000111; // 7: a,b,c ��
            4'd8: LED7S <= 7'b1111111; // 8: ȫ��
            4'd9: LED7S <= 7'b1100111; // 9: a,b,c,f,g ��
			default: LED7S <= 7'b0000000;
        endcase
    end

endmodule