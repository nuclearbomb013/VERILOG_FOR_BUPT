module main(
    input clk_1hz,          // 1Hz ��ʱ�� (����ʱ������)
    input clk_1khz,         // 1000Hz ��Ƶʱ�� (���Ʒ���������)
    input button_1,         // Pulse ��ť - �л�Уʱλ��
    input button_2,         // QD ��ť - ���ӵ�ǰλ��ֵ
    input button_3_raw,     // CLR ��ť (ԭʼ�źţ���Ҫ��ת)
    input switch_clr,       // �ܸ�λ���� (�͵�ƽ��Ч)
    input switch_setting,   // Уʱģʽ����
    input switch_alarm,     // ����ģʽ���� 
    input switch_stopwatch, // ���ģʽ���� 
    input switch_debug1,    // ���Կ���1 - ǿ�Ʒ�������
    input switch_debug2,    // ���Կ���2 (Ԥ��)
    input switch_debug3,    // ���Կ���3 (Ԥ��)
    output [6:0] LED7S_out, 
    output [3:0] LED7S2_out,
    output [3:0] LED7S3_out,
    output [3:0] LED7S4_out,
    output [3:0] LED7S5_out,
    output [3:0] LED7S6_out,
    output beep             // ���������
);
    assign button_3 = ~button_3_raw; // ��ת

    // ��Ƶ���ͽ���������
    // �� 1kHz ʱ�ӷ�Ƶ����
    // - clk_4hz: 4Hz �źţ�������˸��ʾ
    // - rhythm: �����������ź� (ÿ��3��"������")

    reg [9:0] cnt1000;  // 0~999 ���������
    reg clk_4hz;        // 4Hz ������������˸Ч��
    reg rhythm;         // ����������

    always @(posedge clk_1khz or negedge switch_clr) begin
        if (!switch_clr) begin
            cnt1000 <= 10'd0;
        end
        else begin        
            // ���������:0->999->0ѭ��
            if (cnt1000 >= 10'd999) 
                cnt1000 <= 10'd0;
            else 
                cnt1000 <= cnt1000 + 1'b1;

            // 4Hz ��Ƶ: ÿ 250ms ��תһ�� 
            if (cnt1000 == 10'd249 || cnt1000 == 10'd499 || cnt1000 == 10'd749 || cnt1000 == 10'd999)
                clk_4hz <= ~clk_4hz;

            // ����������: ÿ��3����ÿ��100ms
            // 0-100ms: ��, 100-200ms: ͣ, 200-300ms: ��, ...
            if (cnt1000 == 10'd0 || cnt1000 == 10'd200 || cnt1000 == 10'd400)
                rhythm <= 1'b1;
            
            if (cnt1000 == 10'd100 || cnt1000 == 10'd300 || cnt1000 == 10'd500)
                rhythm <= 1'b0;
        end
    end

    // ģʽѡ���߼�
    // ���ȼ�: ��� > ���� > Уʱ > ������
    // mode = 0: ������ģʽ (������ʾʱ��)
    // mode = 1: Уʱģʽ (�ɵ���ʱ��)
    // mode = 2: ����ģʽ (Ԥ��)
    // mode = 3: ���ģʽ (Ԥ��)
    
    wire [1:0] mode;
    assign mode = switch_stopwatch ? 2'd3 :
                  switch_alarm     ? 2'd2 :
                  switch_setting   ? 2'd1 : 2'd0;       


    // �������߼�
    reg [3:0] clock_sec_l;  
    reg [2:0] clock_sec_h;  
    reg [3:0] clock_min_l;
    reg [2:0] clock_min_h; 
    reg [3:0] clock_hour_l;
    reg [1:0] clock_hour_h;

    // ��λʹ���ź�
    wire en_clock_sec_h,en_clock_min_l,en_clock_min_h,en_clock_hour_l,hour_reset;
    
    assign en_clock_sec_h  = (clock_sec_l == 4'd9);                         // ���λ=9ʱ��λ
    assign en_clock_min_l  = (clock_sec_h == 3'd5) && en_clock_sec_h;       // 59��ʱ��λ
    assign en_clock_min_h  = (clock_min_l == 4'd9) && en_clock_min_l;       // X9:59ʱ��λ
    assign en_clock_hour_l = (clock_min_h == 3'd5) && en_clock_min_h;       // 59:59ʱ��λ

    assign hour_reset = (clock_hour_h == 2'd2) && (clock_hour_l == 4'd3); // 23ʱ��λ

    // ʱ�������߼� 
    always @(posedge clk_1hz or negedge switch_clr) begin
        if (!switch_clr) 
            clock_sec_l <= 4'd0;
        else if (load_from_setting) 
            clock_sec_l <= setting_sec_l;
        else case (clock_sec_l)
            4'd9:    clock_sec_l <= 4'd0;
            default: clock_sec_l <= clock_sec_l + 1'b1;
        endcase
    end

    always @(posedge clk_1hz or negedge switch_clr) begin
        if (!switch_clr) 
            clock_sec_h <= 3'd0;
        else if (load_from_setting) 
            clock_sec_h <= setting_sec_h;
        else if (en_clock_sec_h) case (clock_sec_h)
            3'd5:    clock_sec_h <= 3'd0;
            default: clock_sec_h <= clock_sec_h + 1'b1;
        endcase
    end

    always @(posedge clk_1hz or negedge switch_clr) begin
        if (!switch_clr) 
            clock_min_l <= 4'd0;
        else if (load_from_setting) 
            clock_min_l <= setting_min_l;
        else if (en_clock_min_l) case (clock_min_l)
            4'd9:    clock_min_l <= 4'd0;
            default: clock_min_l <= clock_min_l + 1'b1;
        endcase
    end

    always @(posedge clk_1hz or negedge switch_clr) begin
        if (!switch_clr) 
            clock_min_h <= 3'd0;
        else if (load_from_setting) 
            clock_min_h <= setting_min_h;
        else if (en_clock_min_h) case (clock_min_h)
            3'd5:    clock_min_h <= 3'd0;
            default: clock_min_h <= clock_min_h + 1'b1;
        endcase
    end

    always @(posedge clk_1hz or negedge switch_clr) begin
        if (!switch_clr) 
            clock_hour_l <= 4'd0;
        else if (load_from_setting) 
            clock_hour_l <= setting_hour_l;
        else if (en_clock_hour_l) case (1'b1) 
            hour_reset:            clock_hour_l <= 4'd0; 
            (clock_hour_l == 4'd9): clock_hour_l <= 4'd0;
            default:               clock_hour_l <= clock_hour_l + 1'b1;
        endcase
    end

    always @(posedge clk_1hz or negedge switch_clr) begin
        if (!switch_clr) 
            clock_hour_h <= 2'd0;
        else if (load_from_setting) 
            clock_hour_h <= setting_hour_h;
        else if (en_clock_hour_l) case (1'b1)
            hour_reset:            clock_hour_h <= 2'd0;
            (clock_hour_l == 4'd9): clock_hour_h <= clock_hour_h + 1'b1;
            default:               clock_hour_h <= clock_hour_h;
        endcase
    end

    // Уʱ�߼�
    // ��Уʱģʽ�£�����ͨ����ť����ʱ��
    // button_1: �л�����λ�� (�ֵ�->�ָ�->ʱ��->ʱ��)
    // button_2: ���ӵ�ǰλ��ֵ
    // �˳�Уʱģʽʱ�����趨ʱ��ͬ������ʱ��

    reg [3:0] setting_sec_l;
    reg [2:0] setting_sec_h;
    reg [3:0] setting_min_l;
    reg [2:0] setting_min_h;
    reg [3:0] setting_hour_l;
    reg [1:0] setting_hour_h;
    reg [1:0] position;         // ��ǰ����λ�� (0:�ֵ�, 1:�ָ�, 2:ʱ��, 3:ʱ��)
    reg switch_setting_prev;    // Уʱ����ǰһ״̬ (���ڱ��ؼ��)

    // ���Уʱ���ص��½���
    always @(posedge clk_1hz) begin
        switch_setting_prev <= switch_setting;
    end

    // ͬ���ź�: �˳�Уʱģʽʱ����
    wire load_from_setting;
    assign load_from_setting = !switch_setting && switch_setting_prev;

    // �л�����λ�� (����button_1)
    always @(posedge button_1) begin
        if (button_1)
            position <= position + 1;
    end
        
    // ���ӵ�ǰλ��ֵ (����button_2)
    always @(posedge button_2) begin
        if (button_2) begin
            if (mode == 2'd1) begin
                case (position) 
                    // �ֵ�λ: 0-9 ѭ��
                    2'd0: setting_min_l <= (setting_min_l == 4'd9) ? 4'd0 : setting_min_l + 1'b1;
                    // �ָ�λ: 0-5 ѭ��
                    2'd1: setting_min_h <= (setting_min_h == 3'd5) ? 3'd0 : setting_min_h + 1'b1;
                    // ʱ��λ: �迼��24Сʱ����
                    2'd2: begin
                        if (setting_hour_h == 2'd2)
                            // 20-23ʱ��ʱ��λֻ����0-3
                            setting_hour_l <= (setting_hour_l == 4'd3) ? 4'd0 : setting_hour_l + 1'b1;
                        else
                            // 0x-19ʱ��ʱ��λ��0-9
                            setting_hour_l <= (setting_hour_l == 4'd9) ? 4'd0 : setting_hour_l + 1'b1;
                    end
                    
                    // ʱ��λ: 0-2 ѭ�������Զ�����ʱ��λ
                    2'd3: begin
                        // ����������2xʱ����ʱ��λ>3��������Ϊ0
                        if (setting_hour_h == 2'd1 && setting_hour_l > 4'd3)
                            setting_hour_l <= 4'd0;
                        setting_hour_h <= (setting_hour_h == 2'd2) ? 2'd0 : setting_hour_h + 1'b1;
                    end
            endcase
            end
        end
    end 

    // ��ʾ��������
    // ���ݵ�ǰģʽѡ����ʾ����
    // ��Уʱģʽ�£���ǰ����λ����˸ (4Hz)

    wire [3:0] display_1;   // ���λ��ʾֵ
    wire [3:0] display_2;   // ���λ��ʾֵ
    wire [3:0] display_3;   // �ֵ�λ��ʾֵ
    wire [3:0] display_4;   // �ָ�λ��ʾֵ
    wire [3:0] display_5;   // ʱ��λ��ʾֵ
    wire [3:0] display_6;   // ʱ��λ��ʾֵ

    // ����ģʽѡ����ʾԴ: ������ģʽ��ʾclock_*, Уʱģʽ��ʾsetting_*
    assign display_1 = (mode == 2'd0) ? clock_sec_l  : setting_sec_l;
    assign display_2 = (mode == 2'd0) ? {1'b0, clock_sec_h}  : {1'b0, setting_sec_h};
    assign display_3 = (mode == 2'd0) ? clock_min_l  : setting_min_l;
    assign display_4 = (mode == 2'd0) ? {1'b0, clock_min_h}  : {1'b0, setting_min_h};
    assign display_5 = (mode == 2'd0) ? clock_hour_l : setting_hour_l;
    assign display_6 = (mode == 2'd0) ? {2'b00, clock_hour_h} : {2'b00, setting_hour_h};

    // ��˸����: 1��ʾ��λ��Ҫ��˸
    reg [0:5] flicker_mask;

    // LED���: ��˸ʱ��clk_4hz�͵�ƽ�ڼ���ʾ0xF(Ϩ��)
    assign LED7S2_out = ~flicker_mask[1] | clk_4hz ? display_2 : 4'hf;
    assign LED7S3_out = ~flicker_mask[2] | clk_4hz ? display_3 : 4'hf;
    assign LED7S4_out = ~flicker_mask[3] | clk_4hz ? display_4 : 4'hf;
    assign LED7S5_out = ~flicker_mask[4] | clk_4hz ? display_5 : 4'hf;
    assign LED7S6_out = ~flicker_mask[5] | clk_4hz ? display_6 : 4'hf;
    
    // ���λ��Ҫ�߶����� (����λ���ⲿ����������)
    assign LED7S_out = (~flicker_mask[0] | clk_4hz) ? 
        ((display_1 == 4'h0) ? 7'b0111111 :  // 0
         (display_1 == 4'h1) ? 7'b0000110 :  // 1
         (display_1 == 4'h2) ? 7'b1011011 :  // 2
         (display_1 == 4'h3) ? 7'b1001111 :  // 3
         (display_1 == 4'h4) ? 7'b1100110 :  // 4
         (display_1 == 4'h5) ? 7'b1101101 :  // 5
         (display_1 == 4'h6) ? 7'b1111100 :  // 6
         (display_1 == 4'h7) ? 7'b0000111 :  // 7
         (display_1 == 4'h8) ? 7'b1111111 :  // 8
         (display_1 == 4'h9) ? 7'b1100111 :  // 9
         7'b0000000) : 7'b0000000;           // Ϩ��

    // ����Уʱλ��������˸����
    always @(*) begin
        if (mode == 2'd1) begin
            case (position)
                2'd0: flicker_mask = 6'b001000;  // �ֵ�λ��˸
                2'd1: flicker_mask = 6'b000100;  // �ָ�λ��˸
                2'd2: flicker_mask = 6'b000010;  // ʱ��λ��˸
                2'd3: flicker_mask = 6'b000001;  // ʱ��λ��˸
                default: flicker_mask = 6'b000000;
            endcase
        end else begin
            flicker_mask = 6'b000000;  // ��Уʱģʽ����˸
        end
    end


    // �����������߼�
    // ���㱨ʱ: ÿСʱ������5�� (�����ֽ���)
    // ����ģʽ: switch_debug1 ����ʱǿ����

    reg [3:0] beep_timer;   // ��ʱ����ʱ (��λ:��)
    wire beep_enable;       // ������ʹ���ź�
    
    assign beep_enable = (beep_timer != 4'd0) || switch_debug1;
    assign beep = beep_enable && rhythm && clk_1khz;

    always @(posedge clk_1hz) begin
        if (beep_timer > 0) beep_timer <= beep_timer - 1;

        if (en_clock_min_l)
            beep_timer <= 4'd5;
    end


endmodule