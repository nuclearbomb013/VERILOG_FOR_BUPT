module test(
    input clk,
    input clr,          // �ٶ�Ϊ�͵�ƽ��Ч (����ԭ���� negedge)
    output reg [6:0] LED7S,  // ����Ϊ��׼ [6:0] ��ʽ����λ�루�ֶ����룩
    output reg [3:0] LED7S2, // ʮλ�루BCD��
    output reg [3:0] LED7S3, // ��λ�֣�BCD��
    output reg [3:0] LED7S4, // ʮλ�֣�BCD��
    output reg [3:0] LED7S5, // ��λʱ��BCD��
    output reg [3:0] LED7S6  // ʮλʱ��BCD��
);

    reg [5:0] sec;
    reg [5:0] min;
    reg [4:0] hour;
    
    // ���ڸ����������ʱ����
    reg [3:0] sec_unit_val; 

    // ==========================================
    // 1. ʱ�Ӽ����븴λ�߼� (Clock and Reset)
    // ==========================================
    always @(posedge clk or negedge clr) begin
        if (!clr) begin
            // �첽��λ�����¸�λ��ʱ����
            sec <= 0;
            min <= 0;
            hour <= 0;
        end
        else begin
            // ���������߼�
            if (sec >= 59) begin
                sec <= 0;
                if (min >= 59) begin
                    min <= 0;
                    if (hour >= 23)
                        hour <= 0;
                    else
                        hour <= hour + 1;
                end
                else begin
                    min <= min + 1;
                end
            end
            else begin
                sec <= sec + 1;
            end
        end
    end

    // ==========================================
    // 2. ��λ����������߼� (Output Process)
    // ==========================================
    always @(*) begin
        // --- ��λ���벿�� (����������1) ---
        
        // �� (sec)
        sec_unit_val = sec % 10;     // ȡģ�ø�λ
        LED7S2       = sec / 10;     // ������ʮλ
        
        // �� (min)
        LED7S3       = min % 10;     // ��λ
        LED7S4       = min / 10;     // ʮλ
        
        // ʱ (hour)
        LED7S5       = hour % 10;    // ��λ
        LED7S6       = hour / 10;    // ʮλ

        // --- �ֶ����벿�� (�����ĸ�λ) ---
        // �����ǹ��������ǹ�����ȡ����Ӳ���������������ṩ�ı���
        // 4'b0000 -> 7'b1111110 (0x7E, �������������ĸߵ�ƽ�����������ǹ������ĵ͵�ƽ��Ч)
        case (sec_unit_val)
			4'b0000: LED7S <= 7'b1111110; // X"3F"
			4'b0001: LED7S <= 7'b0110000; // X"06"
			4'b0010: LED7S <= 7'b1101101; // X"5B"
			4'b0011: LED7S <= 7'b1111001; // X"4F"
			4'b0100: LED7S <= 7'b0110011; // X"66"
			4'b0101: LED7S <= 7'b1011011; // X"6D"
			4'b0110: LED7S <= 7'b1011111; // X"7D"
			4'b0111: LED7S <= 7'b1110000; // X"07"
			4'b1000: LED7S <= 7'b1111111; // X"7F"
			4'b1001: LED7S <= 7'b1111011; // X"6F"
			default: LED7S <= 7'b0000000;
        endcase
    end

endmodule