module main(
    input clk_1hz,       // 1Hz ��ʱ�� (������ʱ��)
    input clk_1khz,      // 1000Hz ��Ƶʱ�� (���������ֵĽ���)
    input btn_1,     // Pulse 
    input btn_2,     // QD
    input btn_3_raw,     // CLR(��Ҫ��ת)
    input emergncy_stop, // ��ͣ����
    input switch_clr,      // ��λ����
    input simu_hopper_stop, // ©��ֹͣ�ź�
    input simu_hopper_add,  // ©���ֶ�����
    input simu_conveyor_stop, // ���ʹ�ֹͣ�ź�
    input debug_1,
    input debug_2,
    input debug_3,
    input debug_4,
    output [6:0] LED7S_out,
    output [3:0] LED7S2_out,
    output [3:0] LED7S3_out,
    output [3:0] LED7S4_out,
    output [3:0] LED7S5_out,
    output [3:0] LED7S6_out,
    output beep
);

    assign btn_3 = ~btn_3_raw;
    assign hopper_level = ((simu_hopper_stop & state == RUNNING) ? 1'b0 : clk_1hz) | simu_hopper_add; 
    // ©��װҩԭ�źţ�����ÿ���Զ�װҩֻ������״̬����Ч
    wire hopper_signal;
    assign conveyor_signal = ~simu_conveyor_stop; // ���ʹ����������ź�

    // ==========================================
    // ©������ת��
    // ==========================================
    reg hopper_level_prev; // ©��װҩ�ź�
    assign hopper_signal = (hopper_level_prev == 1'b0 && hopper_level == 1'b1);

    always @(posedge clk_1khz) begin
        hopper_level_prev <= hopper_level;
    end

    // ==========================================
    // ��Ƶ
    // ==========================================
    reg [9:0] cnt1k;
    reg clk_4hz; // 4Hz ʱ�ӣ���������ܶ������������˸�ͷ�����
    reg clk_2hz; // 2Hz ʱ�ӣ���������ܷ�����
    reg clk_timer; // ��ʱ��ʱ�ӣ������л���ʱ����©����ʱ��

    always @(posedge clk_1khz) begin
        if (cnt1k == 1000-1) begin
            cnt1k <= 0;
            clk_timer <= ~clk_timer;
        end else
            cnt1k <= cnt1k + 1;
        
        if (cnt1k == 0 || cnt1k == 500)
            clk_2hz <= ~clk_2hz;
        
        if (cnt1k == 0 || cnt1k == 250 || cnt1k == 500 || cnt1k == 750)
            clk_4hz <= ~clk_4hz;
    end

    // ==========================================
    // ��״̬��
    // ==========================================
    
    reg [3:0] target_pills1; // �趨ÿƿҩƬ�� 0~999 ��λ
    reg [3:0] target_pills2; // �趨ÿƿҩƬ�� 0~999 ʮλ
    reg [3:0] target_pills3; // �趨ÿƿҩƬ�� 0~999 ��λ
    reg [3:0] target_bottles1; // �趨��ƿ�� 0~99 ��λ
    reg [3:0] target_bottles2; // �趨��ƿ�� 0~99 ʮλ
    reg [2:0] position; //��λ

    reg [3:0] now_pills1; // ��ǰƿҩƬ�� 0~999 ��λ
    reg [3:0] now_pills2; // ��ǰƿҩƬ�� 0~999 ʮλ
    reg [3:0] now_pills3; // ��ǰƿҩƬ�� 0~999 ��λ
    reg [3:0] now_bottles1; // �Ѿ���ɵ�ƿ�� 0~99 ��λ
    reg [3:0] now_bottles2; // �Ѿ���ɵ�ƿ�� 0~99 ʮλ

    reg [3:0] switch_timer; // �л���ʱ���������ж���һƿ�Ƿ�λ
    wire switch_timer_set; // �л���ʱ�������ź�
    reg [3:0] hopper_timer; // ©����ʱ���������ж�©���Ƿ�ȱ��
    wire hopper_timer_set; // ©����ʱ�������ź�

    parameter [2:0]
        SETTING  = 3'b000, // 0
        RUNNING  = 3'b001, // 1
        SWITCHING = 3'b010, // 2
        DONE     = 3'b011, // 3
        ERROR    = 3'b100, // 4
        FATAL    = 3'b101; // 5
    reg [2:0] state; // ״̬��״̬ 
    reg [2:0] state_next; // ״̬����һ״̬

    always @(posedge clk_1khz or negedge switch_clr) begin
        if (!switch_clr)
            position <= 3'd0;
        else if (btn_1)
            position <= position + 1;
    end

    // ����߼������ж�
    always @(*) begin
        state_next = state;
        if (emergncy_stop) begin
            state_next = FATAL; // ��ͣ���ش����������ش���
        end else begin
            case (state) // ״̬ת������
                SETTING: begin
                    
                end
                RUNNING: begin
                    if (now_pills == target_pills) begin
                        if (now_bottles == target_bottles)
                            state_next = DONE; //װƿ���
                        else 
                            state_next = SWITCHING; //�л�ƿ
                    end else if (hopper_timer == 0) begin
                        state_next = ERROR; // δ�յ�©���źţ���ȱ�ϴ���
                    end
                end
                SWITCHING: begin
                    if (switch_timer == 0) begin
                        if (conveyor_signal)
                            state_next = RUNNING; // ���ʹ��������У���ʼװƿ
                        else
                            state_next = ERROR; // ���ʹ�ֹͣ�������ʹ�����
                    end
                end
                DONE: begin
                    if () // �������ⰴť�ź�
                        state_next = SETTING; // ��λ
                end
                ERROR: begin
                    if (conveyor_signal || hopper_timer != 0) // ���ָ�����
                        state_next = RUNNING; // ��������
                end
                FATAL: begin
                    if () // �������ⰴť�ź�
                        state_next = SETTING; // ��λ
                end
            endcase
        end
    end

    // ʱ���߼�����ת��
    always @(posedge clk_1khz) begin
        if (clk_1khz) begin
            if (state == state_next) begin  
                case (state) // �����߼�
                    SETTING: begin
                        if (btn_3)
                            state_next = RUNNING;
                    end
                    RUNNING: begin
                        // ���м���
                    end
                    SWITCHING: begin
                    end
                    DONE: begin
                    end
                    ERROR: begin
                    end
                    FATAL: begin
                    end
                endcase
            end else begin 
                case (state_next) // ״̬ת��
                    SETTING: begin
                    end
                    RUNNING: begin
                        // ��������̬�����������㣬����������
                    end
                    SWITCHING: begin
                        // �����л�̬�������л���ʱ��2s
                    end
                    DONE: begin
                        
                    end
                    ERROR: begin
                    end
                    FATAL: begin
                    end
                endcase
                state <= state_next;
            end
        end 
    end

    // �л���ʱ���߼�
    always @(posedge clk_timer) begin
        if (switch_timer_set)
            switch_timer <= 2;
        else if (switch_timer != 0)
            switch_timer <= switch_timer - 1;
    end

    // ©����ʱ���߼�
    always @(posedge clk_timer) begin
        if (hopper_timer_set)
            hopper_timer <= 5;
        if (hopper_timer != 0)
            hopper_timer <= hopper_timer - 1;
    end

    // ==========================================
    // SETTING�߼�
    // ==========================================

    // �����߼�
    always @(posedge clk_1khz or negedge switch_clr) begin
    // 1. ��λ��֧�����ȼ���ߣ������κ�״̬����λ�����㣩
        if (!switch_clr) begin
            target_pills1 <= 4'd0;
            target_pills2 <= 4'd0;
            target_pills3 <= 4'd0;
            target_bottles1 <= 4'd0;
            target_bottles2 <= 4'd0;
        end
        // 2. �Ǹ�λ��֧������state==SETTINGʱ����ִ����λ����
        else begin
            // �����޸ģ�����state==SETTING�������ж�
            if (state == SETTING) begin // ֻ���趨״̬�£������������λ
                case (position) 
                    3'd0: target_pills1 <= (target_pills1 == 4'd9) ? 4'd0 : target_pills1 + 1'b1;
                    3'd1: target_pills2 <= (target_pills2 == 4'd9) ? 4'd0 : target_pills2 + 1'b1;
                    3'd2: target_pills3 <= (target_pills3 == 4'd9) ? 4'd0 : target_pills3 + 1'b1; // ������ԭ����
                    3'd3: target_bottles1 <= (target_bottles1 == 4'd9) ? 4'd0 : target_bottles1 + 1'b1; // ������ԭ����
                    3'd4: target_bottles2 <= (target_bottles2 == 4'd9) ? 4'd0 : target_bottles2 + 1'b1;
                endcase

                // ������д��λ�߼�
            end
            // ��SETTING״̬����ִ���κβ���������ԭ��ֵ��VerilogĬ����Ϊ�����������룩
        end
    end

    
    // ==========================================
    // ��ʾ����
    // ==========================================
    // �޸� display_1 ~ display_6 ��ֵ�����޸���ʾ����
    // �޸� flicker_mask[0...5] ��ֵ��������/�ر���˸


    wire [3:0] display_1;
    wire [3:0] display_2;
    wire [3:0] display_3;
    wire [3:0] display_4;
    wire [3:0] display_5;
    wire [3:0] display_6;

    // ������ʾ
    assign display_1 = state;
    assign display_2 = state == SETTING ? target_pills1 : now_pills1;
    assign display_3 = state == SETTING ? target_pills2 : now_pills2;
    assign display_4 = state == SETTING ? target_pills3 : now_pills3;
    assign display_5 = state == SETTING ? target_bottles1 : now_bottles1;
    assign display_6 = state == SETTING ? target_bottles2 : now_bottles2;

    reg [0:5] flicker_mask;

    assign LED7S2_out = ~ flicker_mask[1] | clk_4hz ? display_2 : 4'hf;
    assign LED7S3_out = ~ flicker_mask[2] | clk_4hz ? display_3 : 4'hf;
    assign LED7S4_out = ~ flicker_mask[3] | clk_4hz ? display_4 : 4'hf;
    assign LED7S5_out = ~ flicker_mask[4] | clk_4hz ? display_5 : 4'hf;
    assign LED7S6_out = ~ flicker_mask[5] | clk_4hz ? display_6 : 4'hf;
    assign LED7S_out = (~ flicker_mask[0] | clk_4hz) ?
                        ((display_1 == 0) ? 7'b1001001 : 
                         (display_1 == 1) ? ((anim == 1) ? 7'b0001001 :
                                           (anim == 2) ? 7'b0010010 : 7'b0100100) :
                         (display_1 == 2) ? ((anim == 1) ? 7'b0110000 :
                                           (anim == 2) ? 7'b1000000 : 7'b0000110) :
                         (display_1 == 3) ? ((anim == 1) ? 7'b0111111 :
                                           (anim == 2) ? 7'b0111111 : 7'b0000000) :
                         (display_1 == 4) ? 7'b1111001 :
                         (display_1 == 5) ? 7'b1110001 : 7'b0000000) : 7'b0000000;

    reg [1:0] anim; // 3֡������ʾ

    always @(*) begin
        if(state == SETTING) begin
            case(position)
                3'd0:flicker_mask=6'b010000;
                3'd1:flicker_mask=6'b001000;
                3'd2:flicker_mask=6'b000100;
                3'd3:flicker_mask=6'b000010;
                3'd4:flicker_mask=6'b000001;
                default:flicker_mask=6'b000000;
            endcase
        end else begin
            flicker_mask=6'b000000;
        end
    end

    always @(posedge clk_4hz) begin
        if (anim == 2)
            anim <= 0;
        else
            anim <= anim + 1;
    end


    // ==========================================
    // ����������
    // ==========================================
    reg [4:0] beep_timer; // ��������ʱ��(��λ��250ms)
    assign beep_always = state == DONE;
    assign beep_2hz = state == ERROR;
    assign beep_4hz = state == FATAL;
    
    always @(clk_4hz) begin
        if (beep_timer != 0)
            beep_timer <= beep_timer - 1;
    end

    assign beep = ((beep_timer | beep_always) | (beep_2hz & clk_2hz) | (beep_4hz & clk_4hz)) & clk_1khz;

endmodule

