module test(
    input clk,            // 1Hz ��ʱ�� (������ʱ��)
    input clk_audio,      // 1000Hz ��Ƶʱ�� (���������ֵĽ���)
    input clr,            // ��λ�ź�
    output reg [6:0] LED7S,
    output [3:0] LED7S2,
    output [3:0] LED7S3,
    output [3:0] LED7S4,
    output [3:0] LED7S5,
    output [3:0] LED7S6,
    output beep
);

    // ==========================================
    // 1. ����ʱ��Ĵ���
    // ==========================================
    reg [3:0] sec_l;
    reg [2:0] sec_h;
    reg [3:0] min_l;
    reg [2:0] min_h;
    reg [3:0] hour_l;
    reg [1:0] hour_h;
    
    // ������ʱ�� (���ڿ���ǰ������ж�)
    reg [2:0] start_cnt; 

    // �˿�����
    assign LED7S2 = {1'b0, sec_h};
    assign LED7S3 = min_l;
    assign LED7S4 = {1'b0, min_h};
    assign LED7S5 = hour_l;
    assign LED7S6 = {2'b00, hour_h};

    // ==========================================
    // 2. ������ʹ���߼� (��λ��)
    // ==========================================
    wire en_sec_h, en_min_l, en_min_h, en_hour_l;
    
    assign en_sec_h  = (sec_l == 4'd9);
    assign en_min_l  = (sec_h == 3'd5) && en_sec_h;
    assign en_min_h  = (min_l == 4'd9) && en_min_l;
    assign en_hour_l = (min_h == 3'd5) && en_min_h;
    
    wire hour_reset; 
    assign hour_reset = (hour_h == 2'd2 && hour_l == 4'd3);

    // ==========================================
    // 3. ʱ�������߼� (���ֲ���)
    // ==========================================
    always @(posedge clk or negedge clr) begin
        if (!clr) sec_l <= 4'd0;
        else case (sec_l)
            4'd9:    sec_l <= 4'd0;
            default: sec_l <= sec_l + 1'b1;
        endcase
    end

    always @(posedge clk or negedge clr) begin
        if (!clr) sec_h <= 3'd0;
        else if (en_sec_h) case (sec_h)
            3'd5:    sec_h <= 3'd0;
            default: sec_h <= sec_h + 1'b1;
        endcase
    end

    always @(posedge clk or negedge clr) begin
        if (!clr) min_l <= 4'd0;
        else if (en_min_l) case (min_l)
            4'd9:    min_l <= 4'd0;
            default: min_l <= min_l + 1'b1;
        endcase
    end

    always @(posedge clk or negedge clr) begin
        if (!clr) min_h <= 3'd0;
        else if (en_min_h) case (min_h)
            3'd5:    min_h <= 3'd0;
            default: min_h <= min_h + 1'b1;
        endcase
    end

    always @(posedge clk or negedge clr) begin
        if (!clr) hour_l <= 4'd0;
        else if (en_hour_l) case (1'b1) 
            hour_reset:       hour_l <= 4'd0;
            (hour_l == 4'd9): hour_l <= 4'd0;
            default:          hour_l <= hour_l + 1'b1;
        endcase
    end

    always @(posedge clk or negedge clr) begin
        if (!clr) hour_h <= 2'd0;
        else if (en_hour_l) case (1'b1)
            hour_reset:       hour_h <= 2'd0;
            (hour_l == 4'd9): hour_h <= hour_h + 1'b1;
            default:          hour_h <= hour_h;
        endcase
    end

    // ���������� (����3��ͣ���㹻���ǿ�����2��)
    always @(posedge clk or negedge clr) begin
        if (!clr) start_cnt <= 3'd0;
        else if (start_cnt < 3'd3) start_cnt <= start_cnt + 1'b1;
    end

    // ==========================================
    // 4. ��ʾ���� (���ֲ���)
    // ==========================================
    always @(*) begin
        case (sec_l)
            4'h0: LED7S = 7'b0111111; 4'h1: LED7S = 7'b0000110;
            4'h2: LED7S = 7'b1011011; 4'h3: LED7S = 7'b1001111;
            4'h4: LED7S = 7'b1100110; 4'h5: LED7S = 7'b1101101;
            4'h6: LED7S = 7'b1111100; 4'h7: LED7S = 7'b0000111;
            4'h8: LED7S = 7'b1111111; 4'h9: LED7S = 7'b1100111;
            default: LED7S = 7'b0000000;
        endcase
    end

    // ==========================================
    // 5. �߼��������߼� (���뼶����)
    // ==========================================

    // [Step A] ���崥�����ڣ�ʲôʱ�������죿
    // ���󣺿���ǰ2�� (0,1) �� ����ǰ2�� (0,1)
    reg beep_window;
    always @(*) begin
        // 1. �����Լ� (start_cnt Ϊ 0 �� 1 ʱ)
        if (start_cnt < 3'd2) 
            beep_window = 1'b1;
            
        // 2. ���㱨ʱ (��=00, ��=00��01, �ҿ����Լ��ѽ���)
        else if (min_h == 0 && min_l == 0 && sec_h == 0 && sec_l <= 1)
            beep_window = 1'b1;
            
        else 
            beep_window = 1'b0;
    end

    // [Step B] ��������� (�� 1000Hz ��Ƶʱ������)
    // 0~999 ѭ�������������з�ÿһ��
    reg [9:0] ms_cnt; 
    
    always @(posedge clk_audio or negedge clr) begin
        if (!clr) begin
            ms_cnt <= 10'd0;
        end
        else if (beep_window) begin
            // �ڴ������ڣ�0-999 ѭ������
            if (ms_cnt >= 10'd999) 
                ms_cnt <= 10'd0;
            else 
                ms_cnt <= ms_cnt + 1'b1;
        end
        else begin
            // �����⸴λ����֤�´����ʱ���ͷ��ʼ
            ms_cnt <= 10'd0; 
        end
    end

    // [Step C] ���ɡ������֡�����
    // Ƶ�� 1000Hz -> 1������ = 1ms
    // Ŀ�꣺ÿ�� 3 ��
    reg rhythm;
    always @(*) begin
        // ��1��: 0-100ms
        if (ms_cnt < 100) 
            rhythm = 1'b1;
        // ��2��: 200-300ms
        else if (ms_cnt >= 200 && ms_cnt < 300) 
            rhythm = 1'b1;
        // ��3��: 400-500ms
        else if (ms_cnt >= 400 && ms_cnt < 500) 
            rhythm = 1'b1;
        // ʣ��ʱ�� (500-999ms) ����
        else 
            rhythm = 1'b0;
    end

    // [Step D] �������
    // ֻ���� ������ + ����ΪHigh + ��Ƶʱ���� ʱ����
    assign beep = beep_window & rhythm & clk_audio;

endmodule